`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:41:32 06/01/2016 
// Design Name: 
// Module Name:    Decodificador_VGA 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Decodificador_VGA(
    input clk,
    input [7:0] Contador_1,
	 input [7:0] Contador_2,
	 input [7:0] Contador_3,
	 output reg [7:0] VGA_1,
	 output reg [7:0] VGA_2,
	 output reg [7:0] VGA_3
    );
	 
	 
    always @(posedge clk)
	 begin
       case (Contador_1)
          8'd00: VGA_1 = 8'b00000000;
			 8'd01: VGA_1 = 8'b00000001;
			 8'd02: VGA_1 = 8'b00000010;
			 8'd03: VGA_1 = 8'b00000011;
			 8'd04: VGA_1 = 8'b00000100;
			 8'd05: VGA_1 = 8'b00000101;
			 8'd06: VGA_1 = 8'b00000110;
			 8'd07: VGA_1 = 8'b00000111;
			 8'd08: VGA_1 = 8'b00001000;
			 8'd09: VGA_1 = 8'b00001001;
			 8'd010: VGA_1 = 8'b00010000;
			 8'd011: VGA_1 = 8'b00010001; 
			 8'd012: VGA_1 = 8'b00010010; 
			 8'd013: VGA_1 = 8'b00010011; 
			 8'd014: VGA_1 = 8'b00010100; 
			 8'd015: VGA_1 = 8'b00010101; 
			 8'd016: VGA_1 = 8'b00010110; 
			 8'd017: VGA_1 = 8'b00010111; 
			 8'd018: VGA_1 = 8'b00011000; 
			 8'd019: VGA_1 = 8'b00011001; 
			 8'd020: VGA_1 = 8'b00100000;
			 8'd021: VGA_1 = 8'b00100001;
			 8'd022: VGA_1 = 8'b00100010;
			 8'd023: VGA_1 = 8'b00100011;
			 8'd024: VGA_1 = 8'b00100100;
			 8'd025: VGA_1 = 8'b00100101;
			 8'd026: VGA_1 = 8'b00100110;
			 8'd027: VGA_1 = 8'b00100111;
			 8'd028: VGA_1 = 8'b00101000;
			 8'd029: VGA_1 = 8'b00101001;
			 8'd030: VGA_1 = 8'b00110000;
			 8'd031: VGA_1 = 8'b00110001;
			 8'd032: VGA_1 = 8'b00110010;
			 8'd033: VGA_1 = 8'b00110011;
			 8'd034: VGA_1 = 8'b00110100;
			 8'd035: VGA_1 = 8'b00110101;
			 8'd036: VGA_1 = 8'b00110110;
			 8'd037: VGA_1 = 8'b00110111;
			 8'd038: VGA_1 = 8'b00111000;
			 8'd039: VGA_1 = 8'b00111001;
			 8'd040: VGA_1 = 8'b01000000;
			 8'd041: VGA_1 = 8'b01000001;
			 8'd042: VGA_1 = 8'b01000010;
			 8'd043: VGA_1 = 8'b01000011;
			 8'd044: VGA_1 = 8'b01000100;
			 8'd045: VGA_1 = 8'b01000101;
			 8'd046: VGA_1 = 8'b01000110;
			 8'd047: VGA_1 = 8'b01000111;
			 8'd048: VGA_1 = 8'b01001000;
			 8'd049: VGA_1 = 8'b01001001;
			 8'd050: VGA_1 = 8'b01010000;
			 8'd051: VGA_1 = 8'b01010001;
			 8'd052: VGA_1 = 8'b01010010;
			 8'd053: VGA_1 = 8'b01010011;
			 8'd054: VGA_1 = 8'b01010100; 
			 8'd055: VGA_1 = 8'b01010101;
			 8'd056: VGA_1 = 8'b01010110;
			 8'd057: VGA_1 = 8'b01010111;
			 8'd058: VGA_1 = 8'b01011000;
			 8'd059: VGA_1 = 8'b01011001;
			 8'd060: VGA_1 = 8'b01100000;
			 8'd061: VGA_1 = 8'b01100001;
			 8'd062: VGA_1 = 8'b01100010;
			 8'd063: VGA_1 = 8'b01100011; 
			 8'd064: VGA_1 = 8'b01100100;
			 8'd065: VGA_1 = 8'b01100101;
			 8'd066: VGA_1 = 8'b01100110;
			 8'd067: VGA_1 = 8'b01100111;
			 8'd068: VGA_1 = 8'b01101000;
			 8'd069: VGA_1 = 8'b01101001;
			 8'd070: VGA_1 = 8'b01110000;
			 8'd071: VGA_1 = 8'b01110001;
			 8'd072: VGA_1 = 8'b01110010; 
			 8'd073: VGA_1 = 8'b01110011;
			 8'd074: VGA_1 = 8'b01110100;
			 8'd075: VGA_1 = 8'b01110101;
			 8'd076: VGA_1 = 8'b01110110;
			 8'd077: VGA_1 = 8'b01110111;
			 8'd078: VGA_1 = 8'b01111000;
			 8'd079: VGA_1 = 8'b01111001;
			 8'd080: VGA_1 = 8'b10000000;
			 8'd081: VGA_1 = 8'b10000001;
			 8'd082: VGA_1 = 8'b10000010;
			 8'd083: VGA_1 = 8'b10000011;
			 8'd084: VGA_1 = 8'b10000100;
			 8'd085: VGA_1 = 8'b10000101;
			 8'd086: VGA_1 = 8'b10000110;
			 8'd087: VGA_1 = 8'b10000111;
			 8'd088: VGA_1 = 8'b10001000;
			 8'd089: VGA_1 = 8'b10001001;
			 8'd090: VGA_1 = 8'b10010000;
			 8'd091: VGA_1 = 8'b10010001;
			 8'd092: VGA_1 = 8'b10010010;
			 8'd093: VGA_1 = 8'b10010011;
			 8'd094: VGA_1 = 8'b10010100;
			 8'd095: VGA_1 = 8'b10010101;
			 8'd096: VGA_1 = 8'b10010110;
			 8'd097: VGA_1 = 8'b10010111;
			 8'd098: VGA_1 = 8'b10011000;
			 8'd099: VGA_1 = 8'b10011001;
			 default: VGA_1 = 8'd0;

        endcase
     end
	  
	 always @(posedge clk)
	 begin
       case (Contador_2)
          8'd00: VGA_2 = 8'b00000000;
			 8'd01: VGA_2 = 8'b00000001;
			 8'd02: VGA_2 = 8'b00000010;
			 8'd03: VGA_2 = 8'b00000011;
			 8'd04: VGA_2 = 8'b00000100;
			 8'd05: VGA_2 = 8'b00000101;
			 8'd06: VGA_2 = 8'b00000110;
			 8'd07: VGA_2 = 8'b00000111;
			 8'd08: VGA_2 = 8'b00001000;
			 8'd09: VGA_2 = 8'b00001001;
			 8'd010: VGA_2 = 8'b00010000;
			 8'd011: VGA_2 = 8'b00010001; 
			 8'd012: VGA_2 = 8'b00010010; 
			 8'd013: VGA_2 = 8'b00010011; 
			 8'd014: VGA_2 = 8'b00010100; 
			 8'd015: VGA_2 = 8'b00010101; 
			 8'd016: VGA_2 = 8'b00010110; 
			 8'd017: VGA_2 = 8'b00010111; 
			 8'd018: VGA_2 = 8'b00011000; 
			 8'd019: VGA_2 = 8'b00011001; 
			 8'd020: VGA_2 = 8'b00100000;
			 8'd021: VGA_2 = 8'b00100001;
			 8'd022: VGA_2 = 8'b00100010;
			 8'd023: VGA_2 = 8'b00100011;
			 8'd024: VGA_2 = 8'b00100100;
			 8'd025: VGA_2 = 8'b00100101;
			 8'd026: VGA_2 = 8'b00100110;
			 8'd027: VGA_2 = 8'b00100111;
			 8'd028: VGA_2 = 8'b00101000;
			 8'd029: VGA_2 = 8'b00101001;
			 8'd030: VGA_2 = 8'b00110000;
			 8'd031: VGA_2 = 8'b00110001;
			 8'd032: VGA_2 = 8'b00110010;
			 8'd033: VGA_2 = 8'b00110011;
			 8'd034: VGA_2 = 8'b00110100;
			 8'd035: VGA_2 = 8'b00110101;
			 8'd036: VGA_2 = 8'b00110110;
			 8'd037: VGA_2 = 8'b00110111;
			 8'd038: VGA_2 = 8'b00111000;
			 8'd039: VGA_2 = 8'b00111001;
			 8'd040: VGA_2 = 8'b01000000;
			 8'd041: VGA_2 = 8'b01000001;
			 8'd042: VGA_2 = 8'b01000010;
			 8'd043: VGA_2 = 8'b01000011;
			 8'd044: VGA_2 = 8'b01000100;
			 8'd045: VGA_2 = 8'b01000101;
			 8'd046: VGA_2 = 8'b01000110;
			 8'd047: VGA_2 = 8'b01000111;
			 8'd048: VGA_2 = 8'b01001000;
			 8'd049: VGA_2 = 8'b01001001;
			 8'd050: VGA_2 = 8'b01010000;
			 8'd051: VGA_2 = 8'b01010001;
			 8'd052: VGA_2 = 8'b01010010;
			 8'd053: VGA_2 = 8'b01010011;
			 8'd054: VGA_2 = 8'b01010100; 
			 8'd055: VGA_2 = 8'b01010101;
			 8'd056: VGA_2 = 8'b01010110;
			 8'd057: VGA_2 = 8'b01010111;
			 8'd058: VGA_2 = 8'b01011000;
			 8'd059: VGA_2 = 8'b01011001;
			 8'd060: VGA_2 = 8'b01100000;
			 8'd061: VGA_2 = 8'b01100001;
			 8'd062: VGA_2 = 8'b01100010;
			 8'd063: VGA_2 = 8'b01100011; 
			 8'd064: VGA_2 = 8'b01100100;
			 8'd065: VGA_2 = 8'b01100101;
			 8'd066: VGA_2 = 8'b01100110;
			 8'd067: VGA_2 = 8'b01100111;
			 8'd068: VGA_2 = 8'b01101000;
			 8'd069: VGA_2 = 8'b01101001;
			 8'd070: VGA_2 = 8'b01110000;
			 8'd071: VGA_2 = 8'b01110001;
			 8'd072: VGA_2 = 8'b01110010; 
			 8'd073: VGA_2 = 8'b01110011;
			 8'd074: VGA_2 = 8'b01110100;
			 8'd075: VGA_2 = 8'b01110101;
			 8'd076: VGA_2 = 8'b01110110;
			 8'd077: VGA_2 = 8'b01110111;
			 8'd078: VGA_2 = 8'b01111000;
			 8'd079: VGA_2 = 8'b01111001;
			 8'd080: VGA_2 = 8'b10000000;
			 8'd081: VGA_2 = 8'b10000001;
			 8'd082: VGA_2 = 8'b10000010;
			 8'd083: VGA_2 = 8'b10000011;
			 8'd084: VGA_2 = 8'b10000100;
			 8'd085: VGA_2 = 8'b10000101;
			 8'd086: VGA_2 = 8'b10000110;
			 8'd087: VGA_2 = 8'b10000111;
			 8'd088: VGA_2 = 8'b10001000;
			 8'd089: VGA_2 = 8'b10001001;
			 8'd090: VGA_2 = 8'b10010000;
			 8'd091: VGA_2 = 8'b10010001;
			 8'd092: VGA_2 = 8'b10010010;
			 8'd093: VGA_2 = 8'b10010011;
			 8'd094: VGA_2 = 8'b10010100;
			 8'd095: VGA_2 = 8'b10010101;
			 8'd096: VGA_2 = 8'b10010110;
			 8'd097: VGA_2 = 8'b10010111;
			 8'd098: VGA_2 = 8'b10011000;
			 8'd099: VGA_2 = 8'b10011001;
			 default: VGA_2 = 8'd0;

        endcase
     end
	  
	 always @(posedge clk)
	 begin
       case (Contador_3)
          8'd00: VGA_3 = 8'b00000000;
			 8'd01: VGA_3 = 8'b00000001;
			 8'd02: VGA_3 = 8'b00000010;
			 8'd03: VGA_3 = 8'b00000011;
			 8'd04: VGA_3 = 8'b00000100;
			 8'd05: VGA_3 = 8'b00000101;
			 8'd06: VGA_3 = 8'b00000110;
			 8'd07: VGA_3 = 8'b00000111;
			 8'd08: VGA_3 = 8'b00001000;
			 8'd09: VGA_3 = 8'b00001001;
			 8'd010: VGA_3 = 8'b00010000;
			 8'd011: VGA_3 = 8'b00010001; 
			 8'd012: VGA_3 = 8'b00010010; 
			 8'd013: VGA_3 = 8'b00010011; 
			 8'd014: VGA_3 = 8'b00010100; 
			 8'd015: VGA_3 = 8'b00010101; 
			 8'd016: VGA_3 = 8'b00010110; 
			 8'd017: VGA_3 = 8'b00010111; 
			 8'd018: VGA_3 = 8'b00011000; 
			 8'd019: VGA_3 = 8'b00011001; 
			 8'd020: VGA_3 = 8'b00100000;
			 8'd021: VGA_3 = 8'b00100001;
			 8'd022: VGA_3 = 8'b00100010;
			 8'd023: VGA_3 = 8'b00100011;
			 8'd024: VGA_3 = 8'b00100100;
			 8'd025: VGA_3 = 8'b00100101;
			 8'd026: VGA_3 = 8'b00100110;
			 8'd027: VGA_3 = 8'b00100111;
			 8'd028: VGA_3 = 8'b00101000;
			 8'd029: VGA_3 = 8'b00101001;
			 8'd030: VGA_3 = 8'b00110000;
			 8'd031: VGA_3 = 8'b00110001;
			 8'd032: VGA_3 = 8'b00110010;
			 8'd033: VGA_3 = 8'b00110011;
			 8'd034: VGA_3 = 8'b00110100;
			 8'd035: VGA_3 = 8'b00110101;
			 8'd036: VGA_3 = 8'b00110110;
			 8'd037: VGA_3 = 8'b00110111;
			 8'd038: VGA_3 = 8'b00111000;
			 8'd039: VGA_3 = 8'b00111001;
			 8'd040: VGA_3 = 8'b01000000;
			 8'd041: VGA_3 = 8'b01000001;
			 8'd042: VGA_3 = 8'b01000010;
			 8'd043: VGA_3 = 8'b01000011;
			 8'd044: VGA_3 = 8'b01000100;
			 8'd045: VGA_3 = 8'b01000101;
			 8'd046: VGA_3 = 8'b01000110;
			 8'd047: VGA_3 = 8'b01000111;
			 8'd048: VGA_3 = 8'b01001000;
			 8'd049: VGA_3 = 8'b01001001;
			 8'd050: VGA_3 = 8'b01010000;
			 8'd051: VGA_3 = 8'b01010001;
			 8'd052: VGA_3 = 8'b01010010;
			 8'd053: VGA_3 = 8'b01010011;
			 8'd054: VGA_3 = 8'b01010100; 
			 8'd055: VGA_3 = 8'b01010101;
			 8'd056: VGA_3 = 8'b01010110;
			 8'd057: VGA_3 = 8'b01010111;
			 8'd058: VGA_3 = 8'b01011000;
			 8'd059: VGA_3 = 8'b01011001;
			 8'd060: VGA_3 = 8'b01100000;
			 8'd061: VGA_3 = 8'b01100001;
			 8'd062: VGA_3 = 8'b01100010;
			 8'd063: VGA_3 = 8'b01100011; 
			 8'd064: VGA_3 = 8'b01100100;
			 8'd065: VGA_3 = 8'b01100101;
			 8'd066: VGA_3 = 8'b01100110;
			 8'd067: VGA_3 = 8'b01100111;
			 8'd068: VGA_3 = 8'b01101000;
			 8'd069: VGA_3 = 8'b01101001;
			 8'd070: VGA_3 = 8'b01110000;
			 8'd071: VGA_3 = 8'b01110001;
			 8'd072: VGA_3 = 8'b01110010; 
			 8'd073: VGA_3 = 8'b01110011;
			 8'd074: VGA_3 = 8'b01110100;
			 8'd075: VGA_3 = 8'b01110101;
			 8'd076: VGA_3 = 8'b01110110;
			 8'd077: VGA_3 = 8'b01110111;
			 8'd078: VGA_3 = 8'b01111000;
			 8'd079: VGA_3 = 8'b01111001;
			 8'd080: VGA_3 = 8'b10000000;
			 8'd081: VGA_3 = 8'b10000001;
			 8'd082: VGA_3 = 8'b10000010;
			 8'd083: VGA_3 = 8'b10000011;
			 8'd084: VGA_3 = 8'b10000100;
			 8'd085: VGA_3 = 8'b10000101;
			 8'd086: VGA_3 = 8'b10000110;
			 8'd087: VGA_3 = 8'b10000111;
			 8'd088: VGA_3 = 8'b10001000;
			 8'd089: VGA_3 = 8'b10001001;
			 8'd090: VGA_3 = 8'b10010000;
			 8'd091: VGA_3 = 8'b10010001;
			 8'd092: VGA_3 = 8'b10010010;
			 8'd093: VGA_3 = 8'b10010011;
			 8'd094: VGA_3 = 8'b10010100;
			 8'd095: VGA_3 = 8'b10010101;
			 8'd096: VGA_3 = 8'b10010110;
			 8'd097: VGA_3 = 8'b10010111;
			 8'd098: VGA_3 = 8'b10011000;
			 8'd099: VGA_3 = 8'b10011001;
			 default: VGA_3 = 8'd0;

        endcase
     end

endmodule
